interface mux_if;
 logic [3:0] i0,i1,i2,i3;
 logic [1:0] sel;
 logic [3:0] y;
endinterface