package mux_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

 `include "trans.sv"

 `include "seq.sv"
 `include "mon.sv"
 `include "drv.sv"
 `include "seqr.sv"

 `include "agt.sv"
 `include "scoreboard.sv"
 `include "env.sv"

 `include "test.sv"

endpackage